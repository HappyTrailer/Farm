    ����          Assembly-CSharp   qSystem.Collections.Generic.List`1[[Item, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  Item[]   	   >   J          �   Item   	   	   	   	   	   		   	
   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	    	!   	"   	#   	$   	%   	&   	'   	(   	)   	*   	+   	,   	-   	.   	/   	0   	1   	2   	3   	4   	5   	6   	7   	8   	9   	:   	;   	<   	=   	>   	?   	@   	A   B   ItemInInventory   item_idid	itemPriceitemNameitemType
spritePath	itemCount              K   B   PotatoC   seadD   plUnicum               2   E   TomatF   harvestG   fruit1
               2   H   Tomat	F   I   fruit1               2   J   Tomat	F   K   fruit1
               2   L   Tomat	F   M   fruit1
   	            2   N   Tomat	F   O   fruit1
   
            2   P   Tomat	F   Q   fruit1
               2   R   Tomat	F   S   fruit1
               2   T   Tomat	F   U   fruit1
         	      2   V   Tomat	F   W   fruit1
         
      2   X   Tomat	F   Y   fruit1
               2   Z   Tomat	F   [   fruit1
               2   \   Tomat	F   ]   fruit1
               2   ^   Tomat	F   _   fruit1
               2   `   Tomat	F   a   fruit1
               2   b   Tomat	F   c   fruit1
               2   d   Tomat	F   e   fruit1
               2   f   Tomat	F   g   fruit1
               2   h   Tomat	F   i   fruit1
               2   j   Tomat	F   k   fruit1
               2   l   Tomat	F   m   fruit1
               2   n   Tomat	F   o   fruit1
               2   p   Tomat	F   q   fruit1
               2   r   Tomat	F   s   fruit1               2   t   Tomat	F   u   fruit1
               2   v   Tomat	F   w   fruit1
               2   x   Tomat	F   y   fruit1
               2   z   Tomat	F   {   fruit1
                2   |   Tomat	F   }   fruit1
   !            2   ~   Tomat	F      fruit1
   "            2   �   Tomat	F   �   fruit1
   #            2   �   Tomat	F   �   fruit1
   $             2   �   Tomat	F   �   fruit1
   %      !      2   �   Tomat	F   �   fruit1
   &      "      2   �   Tomat	F   �   fruit1
   '      #      2   �   Tomat	F   �   fruit1
   (      $      2   �   Tomat	F   �   fruit1
   )      %      2   �   Tomat	F   �   fruit1
   *      &      2   �   Tomat	F   �   fruit1
   +      '      2   �   Tomat	F   �   fruit1
   ,      (      2   �   Tomat	F   �   fruit1
   -      )      2   �   Tomat	F   �   fruit1
   .      *      2   �   Tomat	F   �   fruit1
   /      +      2   �   Tomat	F   �   fruit1
   0      ,      2   �   Tomat	F   �   fruit1   1      -      2   �   Tomat	F   �   fruit1
   2      .      2   �   Tomat	F   �   fruit1
   3      /      2   �   Tomat	F   �   fruit1
   4      0      2   �   Tomat	F   �   fruit1
   5      1      2   �   Tomat	F   �   fruit1
   6      2      2   �   Tomat	F   �   fruit1
   7      3      2   �   Tomat	F   �   fruit1
   8      4      2   �   Tomat	F   �   fruit1
   9      5      2   �   Tomat	F   �   fruit1
   :      6      2   �   Tomat	F   �   fruit1
   ;      7      2   �   Tomat	F   �   fruit1
   <      8      2   �   Tomat	F   �   fruit1
   =      9      2   �   Tomat	F   �   fruit1
   >      :      2   �   Tomat	F   �   fruit1
   ?      ;      2   �   Tomat	F   �   fruit1
   @      <      2   �   Tomat	F   �   fruit1
   A      =      2   �   Tomat	F   �   fruit1
   