    ����          Assembly-CSharp   wSystem.Collections.Generic.List`1[[fildEvents, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  fildEvents[]   	                      
fildEvents   