    ����          Assembly-CSharp   qSystem.Collections.Generic.List`1[[Item, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  Item[]   	                   Item   	   	   

   ItemInInventory   item_idid	itemPriceitemNameitemType
spritePath	itemCount                    Репа   sead	                     	      harvest	      