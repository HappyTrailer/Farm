    ����          Assembly-CSharp   qSystem.Collections.Generic.List`1[[Item, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  Item[]   	                   Item   	   	   	   
   ItemInInventory   id	itemPriceitemNameitemType
spritePath	itemCount         2      Tomat   sead	   pl4            K   
   Potato	      plUnicum            2      Tomat   harvest   fruit12   