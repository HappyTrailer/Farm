    ����          Assembly-CSharp   vSystem.Collections.Generic.List`1[[SaveField, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  SaveField[]   	   2   2          @   	SaveField   	   	   	   	   	   		   	
   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	    	!   	"   	#   	$   	%   	&   	'   	(   	)   	*   	+   	,   	-   	.   	/   	0   	1   	2   	3   	4   	5      	SaveField   idFildlockeddigwateringweed
fertilizerverminsownwateringTime
timeFactorplant          	SavePlant                    A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
	                   A  �?

                   A  �?
                   A  �?
                   A  �?
      	             A  �?
      
             A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                   A  �?
                    A  �?
!                   A  �?
"                   A  �?
#                   A  �?
$                    A  �?
%      !             A  �?
&      "             A  �?
'      #             A  �?
(      $             A  �?
)      %             A  �?
*      &             A  �?
+      '             A  �?
,      (             A  �?
-      )             A  �?
.      *             A  �?
/      +             A  �?
0      ,             A  �?
1      -             A  �?
2      .             A  �?
3      /             A  �?
4      0             A  �?
5      1             A  �?
