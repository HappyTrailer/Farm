    ����          Assembly-CSharp   qSystem.Collections.Generic.List`1[[Item, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  Item[]   	   A   G          �   Item   	   	   	   	   	   		   	
   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	    	!   	"   	#   	$   	%   	&   	'   	(   	)   	*   	+   	,   	-   	.   	/   	0   	1   	2   	3   	4   	5   	6   	7   	8   	9   	:   	;   	<   	=   	>   	?   	@   	A   	B   	C   	D   ?   ItemInInventory   item_idid	itemPriceitemNameitemType
spritePath	itemCount              K   E   PotatoF   seadG   plUnicum               2   H   TomatI   harvestJ   fruit1
               2   K   Tomat	I   L   fruit1
               2   M   Tomat	I   N   fruit1
               2   O   Tomat	I   P   fruit1
   	            2   Q   Tomat	I   R   fruit1
   
            2   S   Tomat	I   T   fruit1
               2   U   Tomat	I   V   fruit1
               2   W   Tomat	I   X   fruit1
         	      2   Y   Tomat	I   Z   fruit1
         
      2   [   Tomat	I   \   fruit1
               2   ]   Tomat	I   ^   fruit1
               2   _   Tomat	I   `   fruit1
               2   a   Tomat	I   b   fruit1
               2   c   Tomat	I   d   fruit1
               2   e   Tomat	I   f   fruit1
               2   g   Tomat	I   h   fruit1
               2   i   Tomat	I   j   fruit1
               2   k   Tomat	I   l   fruit1
               2   m   Tomat	I   n   fruit1
               2   o   Tomat	I   p   fruit1
               2   q   Tomat	I   r   fruit1
               2   s   Tomat	I   t   fruit1
               2   u   Tomat	I   v   fruit1
               2   w   Tomat	I   x   fruit1
               2   y   Tomat	I   z   fruit1
               2   {   Tomat	I   |   fruit1
               2   }   Tomat	I   ~   fruit1
                2      Tomat	I   �   fruit1
   !            2   �   Tomat	I   �   fruit1
   "            2   �   Tomat	I   �   fruit1
   #            2   �   Tomat	I   �   fruit1
   $             2   �   Tomat	I   �   fruit1
   %      !      2   �   Tomat	I   �   fruit1
   &      "      2   �   Tomat	I   �   fruit1
   '      #      2   �   Tomat	I   �   fruit1
   (      $      2   �   Tomat	I   �   fruit1
   )      %      2   �   Tomat	I   �   fruit1
   *      &      2   �   Tomat	I   �   fruit1
   +      '      2   �   Tomat	I   �   fruit1
   ,      (      2   �   Tomat	I   �   fruit1
   -      )      2   �   Tomat	I   �   fruit1
   .      *      2   �   Tomat	I   �   fruit1
   /      +      2   �   Tomat	I   �   fruit1
   0      ,      2   �   Tomat	I   �   fruit1
   1      -      2   �   Tomat	I   �   fruit1
   2      .      2   �   Tomat	I   �   fruit1
   3      /      2   �   Tomat	I   �   fruit1
   4      0      2   �   Tomat	I   �   fruit1
   5      1      2   �   Tomat	I   �   fruit1
   6      2      2   �   Tomat	I   �   fruit1
   7      3      2   �   Tomat	I   �   fruit1
   8      4      2   �   Tomat	I   �   fruit1
   9      5      2   �   Tomat	I   �   fruit1
   :      6      2   �   Tomat	I   �   fruit1
   ;      7      2   �   Tomat	I   �   fruit1
   <      8      2   �   Tomat	I   �   fruit1
   =      9      2   �   Tomat	I   �   fruit1
   >      :      2   �   Tomat	I   �   fruit1
   ?      ;      2   �   Tomat	I   �   fruit1
   @      <      2   �   Tomat	I   �   fruit1
   A      =      2   �   Tomat	I   �   fruit1
   B      >      2   �   Tomat	I   �   fruit1
   C      ?      2   �   Tomat	I   �   fruit1
   D      @      2   �   Tomat	I   �   fruit1   