    ����          Assembly-CSharp   wSystem.Collections.Generic.List`1[[fildEvents, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  fildEvents[]   	                   
fildEvents   	   	   	   	   	      
fildEvents   _fild_time_type        O4�3 0Ԉ	   weed         �u9 0Ԉ
   vermin         �u� 0Ԉ   watering         Sc�� 0Ԉ	             ϶� 0Ԉ	   