    ����          Assembly-CSharp   qSystem.Collections.Generic.List`1[[Item, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  Item[]   	   ;   M          �   Item   	   	   	   	   	   		   	
   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	    	!   	"   	#   	$   	%   	&   	'   	(   	)   	*   	+   	,   	-   	.   	/   	0   	1   	2   	3   	4   	5   	6   	7   	8   	9   	:   	;   	<   	=   	>   E   ItemInInventory   item_idid	itemPriceitemNameitemType
spritePath	itemCount              K   ?   Potato@   seadA   plUnicum               2   B   TomatC   harvestD   fruit1
               2   E   Tomat	C   F   fruit1               2   G   Tomat	C   H   fruit1
               2   I   Tomat	C   J   fruit1
   	            2   K   Tomat	C   L   fruit1
   
            2   M   Tomat	C   N   fruit1
               2   O   Tomat	C   P   fruit1
               2   Q   Tomat	C   R   fruit1
         	      2   S   Tomat	C   T   fruit1
         
      2   U   Tomat	C   V   fruit1
               2   W   Tomat	C   X   fruit1
               2   Y   Tomat	C   Z   fruit1
               2   [   Tomat	C   \   fruit1
               2   ]   Tomat	C   ^   fruit1
               2   _   Tomat	C   `   fruit1
               2   a   Tomat	C   b   fruit1
               2   c   Tomat	C   d   fruit1
               2   e   Tomat	C   f   fruit1
               2   g   Tomat	C   h   fruit1
               2   i   Tomat	C   j   fruit1               2   k   Tomat	C   l   fruit1
               2   m   Tomat	C   n   fruit1
               2   o   Tomat	C   p   fruit1
               2   q   Tomat	C   r   fruit1
               2   s   Tomat	C   t   fruit1
               2   u   Tomat	C   v   fruit1
               2   w   Tomat	C   x   fruit1
                2   y   Tomat	C   z   fruit1
   !            2   {   Tomat	C   |   fruit1
   "             2   }   Tomat	C   ~   fruit1
   #      !      2      Tomat	C   �   fruit1
   $      "      2   �   Tomat	C   �   fruit1
   %      #      2   �   Tomat	C   �   fruit1
   &      $      2   �   Tomat	C   �   fruit1
   '      %      2   �   Tomat	C   �   fruit1
   (      &      2   �   Tomat	C   �   fruit1
   )      '      2   �   Tomat	C   �   fruit1
   *      (      2   �   Tomat	C   �   fruit1
   +      )      2   �   Tomat	C   �   fruit1
   ,      *      2   �   Tomat	C   �   fruit1
   -      +      2   �   Tomat	C   �   fruit1   .      ,      2   �   Tomat	C   �   fruit1	   /      -      2   �   Tomat	C   �   fruit1
   0      .      2   �   Tomat	C   �   fruit1
   1      /      2   �   Tomat	C   �   fruit1
   2      0      2   �   Tomat	C   �   fruit1
   3      1      2   �   Tomat	C   �   fruit1
   4      2      2   �   Tomat	C   �   fruit1
   5      3      2   �   Tomat	C   �   fruit1
   6      4      2   �   Tomat	C   �   fruit1
   7      5      2   �   Tomat	C   �   fruit1
   8      6      2   �   Tomat	C   �   fruit1
   9      7      2   �   Tomat	C   �   fruit1
   :      8      2   �   Tomat	C   �   fruit1
   ;      9      2   �   Tomat	C   �   fruit1
   <      :      2   �   Tomat	C   �   fruit1
   =      ;      2   �   Tomat	C   �   fruit1
   >      <      2   �   Tomat	C   �   fruit1
   