    ����          Assembly-CSharp   qSystem.Collections.Generic.List`1[[Item, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  Item[]   	   I   _          �   Item   	   	   	   	   	   		   	
   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	    	!   	"   	#   	$   	%   	&   	'   	(   	)   	*   	+   	,   	-   	.   	/   	0   	1   	2   	3   	4   	5   	6   	7   	8   	9   	:   	;   	<   	=   	>   	?   	@   	A   	B   	C   	D   	E   	F   	G   	H   	I   	J   	K   	L   7   ItemInInventory   item_idid	itemPriceitemNameitemType
spritePath	itemCount              2   M   TomatN   harvestO   fruit1
               2   P   Tomat	N   Q   fruit1
               2   R   Tomat	N   S   fruit1
               2   T   Tomat	N   U   fruit1
               2   V   Tomat	N   W   fruit1
   	            2   X   Tomat	N   Y   fruit1
   
            2   Z   Tomat	N   [   fruit1
               2   \   Tomat	N   ]   fruit1
               2   ^   Tomat	N   _   fruit1
         	      2   `   Tomat	N   a   fruit1
         
      2   b   Tomat	N   c   fruit1
               2   d   Tomat	N   e   fruit1
               2   f   Tomat	N   g   fruit1
               2   h   Tomat	N   i   fruit1
               2   j   Tomat	N   k   fruit1
               2   l   Tomat	N   m   fruit1
               2   n   Tomat	N   o   fruit1
               2   p   Tomat	N   q   fruit1
               2   r   Tomat	N   s   fruit1
               2   t   Tomat	N   u   fruit1
               2   v   Tomat	N   w   fruit1
               2   x   Tomat	N   y   fruit1
               2   z   Tomat	N   {   fruit1
               2   |   Tomat	N   }   fruit1
               2   ~   Tomat	N      fruit1
               2   �   Tomat	N   �   fruit1
               2   �   Tomat	N   �   fruit1
               2   �   Tomat	N   �   fruit1
                2   �   Tomat	N   �   fruit1
   !            2   �   Tomat	N   �   fruit1
   "            2   �   Tomat	N   �   fruit1
   #            2   �   Tomat	N   �   fruit1
   $             2   �   Tomat	N   �   fruit1
   %      !      2   �   Tomat	N   �   fruit1
   &      "      2   �   Tomat	N   �   fruit1
   '      #      2   �   Tomat	N   �   fruit1
   (      $      2   �   Tomat	N   �   fruit1
   )      %      2   �   Tomat	N   �   fruit1
   *      &      2   �   Tomat	N   �   fruit1
   +      '      2   �   Tomat	N   �   fruit1
   ,      (      2   �   Tomat	N   �   fruit1
   -      )      2   �   Tomat	N   �   fruit1
   .      *      2   �   Tomat	N   �   fruit1
   /      +      2   �   Tomat	N   �   fruit1
   0      ,      2   �   Tomat	N   �   fruit1
   1      -      2   �   Tomat	N   �   fruit1
   2      .      2   �   Tomat	N   �   fruit1
   3      /      2   �   Tomat	N   �   fruit1
   4      0      2   �   Tomat	N   �   fruit1
   5      1      2   �   Tomat	N   �   fruit1
   6      2      2   �   Tomat	N   �   fruit1
   7      3      2   �   Tomat	N   �   fruit1
   8      4      2   �   Tomat	N   �   fruit1
   9      5      2   �   Tomat	N   �   fruit1
   :      6      2   �   Tomat	N   �   fruit1
   ;      7      2   �   Tomat	N   �   fruit1
   <      8      2   �   Tomat	N   �   fruit1
   =      9      2   �   Tomat	N   �   fruit1
   >      :      K   �   Potato�   harvest�   fruit2
   ?      ;      2   �   Tomat�   sead�   pl4   @      <      2   �   Tomat�   harvest�   fruit1
   A      =      2   �   Tomat	�   �   fruit1
   B      >      2   �   Tomat	�   �   fruit1
   C      ?      2   �   Tomat	�   �   fruit1
   D      @      2   �   Tomat	�   �   fruit1
   E      A      2   �   Tomat	�   �   fruit1	   F      B      2   �   Tomat	�   �   fruit1
   G      C      2   �   Tomat	�   �   fruit1
   H      D      2   �   Tomat	�   �   fruit1   I      E      2   �   Tomat	�   �   fruit1
   J      F      2   �   Tomat	�   �   fruit1
   K      G      2   �   Tomat	�   �   fruit1   L      H      K   �   Potato�   harvest�   fruit2   