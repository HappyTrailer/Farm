    ����          Assembly-CSharp   vSystem.Collections.Generic.List`1[[SaveField, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  SaveField[]   	   2   2          @   	SaveField   	   	   	   	   	   		   	
   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	   	    	!   	"   	#   	$   	%   	&   	'   	(   	)   	*   	+   	,   	-   	.   	/   	0   	1   	2   	3   	4   	5      	SaveField   idFildlockeddigwateringweed
fertilizerverminsownwateringTime
timeFactorplant          	SavePlant                  A��L?	6                   A  �?	7                    A��L?	8                     A  �?
                  A  �?
	                  A  �?

                  A  �?
                  A  �?
                  A  �?
      	            A  �?
      
            A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                  A  �?
                   A  �?
!                  A  �?
"                  A  �?
#                  A  �?
$                   A  �?
%      !            A  �?
&      "            A  �?
'      #            A  �?
(      $            A  �?
)      %            A  �?
*      &            A  �?
+      '            A  �?
,      (            A  �?
-      )            A  �?
.      *            A  �?
/      +            A  �?
0      ,            A  �?
1      -            A  �?
2      .            A  �?
3      /            A  �?
4      0            A  �?
5      1            A  �?
6   	SavePlant   fruitIdnameoldTimeFactormincountFruitmaxcountFruititerationFruitcountExpiriensstageOnestageTwo
stageThree	stageFourbuffStageThreebuffStageFourcurrentStageplantedgrowingstage                     9   Репа   ����?             ��A@  @A  @A  @A  pA  pA    :   stage17   6      	9         �?             r�-@  @A  @A  @A  pA  pA    	:   8   6      	9      ����?             �	@  @A  @A  @A  pA  pA    	:   